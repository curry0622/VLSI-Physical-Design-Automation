# Company Name: Silicon Canvas
# Product Name: Laker
# Software Version: 2021.03

VERSION 5.6 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.01 ;

LAYER CONT
  TYPE CUT ;
END CONT

LAYER PO1
  TYPE MASTERSLICE ;
END PO1

LAYER ME1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.72 ;
  WIDTH 0.24 ;
  OFFSET 0 ;
  SPACING 0.24 ;
END ME1

LAYER VI1
  TYPE CUT ;
END VI1

LAYER ME2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.72 ;
  WIDTH 0.28 ;
  OFFSET 0 ;
  SPACING 0.28 ;
END ME2

LAYER VI2
  TYPE CUT ;
END VI2

LAYER ME3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.72 ;
  WIDTH 0.28 ;
  OFFSET 0 ;
  SPACING 0.28 ;
END ME3

LAYER VI3
  TYPE CUT ;
END VI3

LAYER ME4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.72 ;
  WIDTH 0.28 ;
  OFFSET 0 ;
  SPACING 0.28 ;
END ME4

LAYER VI4
  TYPE CUT ;
END VI4

LAYER ME5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.72 ;
  WIDTH 0.28 ;
  OFFSET 0 ;
  SPACING 0.28 ;
END ME5

LAYER VI5
  TYPE CUT ;
END VI5

LAYER ME6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 2.2 ;
  WIDTH 1.2 ;
  OFFSET 0 ;
  SPACING 1 ;
END ME6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

END LIBRARY
