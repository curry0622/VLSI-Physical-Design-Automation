/users/course/2022F/PDA13400000/g111062625/VLSI-PDA-HW-2022/HW1/test4/NangateOpenCellLibrary.lef