/users/course/2022F/PDA13400000/g111062625/VLSI-PDA-HW-2022/HW1/tests/5ns_0.8_high_on/NangateOpenCellLibrary.lef