/users/course/2022F/PDA13400000/g111062625/HW1/NangateOpenCellLibrary.lef